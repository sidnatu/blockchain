module miner_fsm (

input logic clk,
input logic rst,
input logic cmd_valid,

output logic not_found

);











endmodule